// ADS131A0x Driver Development Project
// Interface: 	SPI Protocol, Cyclone 10 LP Intel FPGA
// Author: 		Dennis Wong
// Date:			6/2/2025 


/* Top Module */
module ADS131A0X (
    input 				system_clock, 			// 50 Mhz system clock
	 input				reset_n,					// Reset activated by push button
	 output 				[3:0]led,				// leds 
	 
	 /* SPI  */
	 output 				SPI_MOSI,				// SPI MOSI
	 input 				SPI_MISO,				// SPI MISO
	 output				SPI_CS,					//	SPI CS
	 output 				SPI_SCLK,				// SPI SCLK
	 output 				SPI_RESET,				// SPI_RESET
	 
	 /* SPI Signals */
	input					adc_init,				// Trigger signal to init the adc					- for simulation (consider removing in final design)
	input 				adc_ready,				// Trigger signal to send SPI transaction			- for simulation (consider removing in final design)
	output [2:0]		state,					// Keeps track of the current state of SPI 		- for debugging (remove in final design)
	output 				adc_init_completed_z // Keeps track of the init progress of the ADC 	- for debugging (remove in final design)
);

wire synthesized_clock_1Mhz;					// 1Mhz clock for heartbeat
wire synthesized_clock_4Mhz;					// 4Mhz clock for SPI_Clock
wire spi_sclk;										// SPI Clock

/* Clock Synthesis Instance */
clock_synthesizer clock_synthesizer_uut_1
(
    .input_clock(system_clock), 							// input clock  - 50 Mhz
	 .clock_pol(led[1])										// output clock to led0 @ 1Mhz
);

/* Clock Synthesizer for SPI with CS Consideration */
spi_sclk_generator spi_sclk_generator_uut (
    .clk(system_clock),      // System clock - 50Mhz
    .cs(SPI_CS),       // Chip Select (Active LOW)
    .sclk(led[3])      // SPI Clock output
);

/* Heartbeat Instance */
heartbeat heartbeat_uut(
    .input_clock(system_clock), 							// 50 Mhz system clock
	 .clock_pol(led[0])										// output clock to led0 @ 1Mhz
);


/* SPI_Master Instance */
SPI_Master SPI_Master_uut
(
	.system_clock(system_clock),							// System Clock from FPGA - 50Mhz
	.reset_n(reset_n),										// Reset_n manually activated by push button	
	.SPI_MOSI(SPI_MOSI),										// SPI MOSI
	.SPI_MISO(SPI_MISO),										// SPI MISO
	.SPI_CS(SPI_CS),											//	SPI CS
	.SPI_SCLK(spi_sclk),										// SPI SCLK
	.SPI_RESET(SPI_RESET),
	
	/* Non crucial Signals (for simulation and debugging) */
	.adc_init_completed_z(adc_init_completed_z),
	.state(state),												// Keeps track of the current state of SPI
	.adc_init(adc_init),										// Trigger signal to init the adc
	.adc_ready(adc_ready)									// Trigger signal to send SPI transaction
);

// assign led[3] = 1'b1;										// assign led to low
assign led[2] = spi_sclk;									// assign led[2] to 4.167Mhz (debug)

assign SPI_SCLK = spi_sclk;								// assign the SPI_SCLK to 4.167Mhz generated by SPI_Master module 

endmodule
