// ADS131A0x Driver Development Project
// Interface: 	SPI Protocol, Cyclone 10 LP Intel FPGA
// Author: 		Dennis Wong
// Date:			6/2/2025 


/* Top Module */
module ADS131A0X (
    input 				system_clock, 			// 50 Mhz system clock
	 input				reset_n,					// Reset activated by push button
	 output 				[3:0]led,				// leds 
	 
	 /* SPI  */
	 output 				SPI_MOSI,				// SPI MOSI
	 input 				SPI_MISO,				// SPI MISO
	 output				SPI_CS,					//	SPI CS
	 output 				SPI_SCLK,					// SPI SCLK
	 
	 /* SPI Signals */
	input					adc_init,				// Trigger signal to init the adc
	input 				adc_ready,				// Trigger signal to send SPI transaction
	output [2:0]		state					// Keeps track of the current state of SPI
);

wire synthesized_clock_1Mhz;					// 1Mhz clock for heartbeat
wire synthesized_clock_4Mhz;					// 4Mhz clock for SPI_Clock
wire spi_sclk;										// SPI Clock

/* Clock Synthesis Instance */
clock_synthesizer clock_synthesizer_uut_1
(
    .input_clock(system_clock), 							// input clock  - 50 Mhz
	 .clock_pol(led[1])										// output clock - 1Mhz 
);

/* Heartbeat Instance */
heartbeat heartbeat_uut(
    .input_clock(system_clock), 							// 50 Mhz system clock
	 .clock_pol(led[0])										// leds 
);


/* SPI_Master Instance */
SPI_Master 
(
	.system_clock(system_clock),							// System Clock from FPGA - 50Mhz
	.reset_n(reset_n),										// Reset_n manually activated by push button	
	.adc_init(adc_init),										// Trigger signal to init the adc
	.adc_ready(adc_ready),									// Trigger signal to send SPI transaction
	.state(state),												// Keeps track of the current state of SPI
	
	.SPI_MOSI(SPI_MOSI),										// SPI MOSI
	.SPI_MISO(SPI_MISO),										// SPI MISO
	.SPI_CS(SPI_CS),											//	SPI CS
	.SPI_SCLK(spi_sclk)										// SPI SCLK
);

assign led[3] = 1'b1;										// assign led to low
assign led[2] = spi_sclk;									// assign led[2] to 4.167Mhz (debug)

assign SPI_SCLK = spi_sclk;								// assign the SPI_SCLK to 4.167Mhz generated by SPI_Master module 

endmodule
